-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
configuration descrambler_config of descrambler is
   for struct
   end for;
end descrambler_config;
