-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
configuration channel_selection_config of channel_selection is
   for struct
   end for;
end channel_selection_config;
