configuration ANDgate4_config of ANDgate4 is
   for untitled
   end for;
end ANDgate4_config;