configuration ORgate_config of ORgate is
   for untitled
   end for;
end ORgate_config;