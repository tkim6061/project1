-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
configuration scrambler2_config of scrambler2 is
   for struct
   end for;
end scrambler2_config;
