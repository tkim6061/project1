configuration ANDgate5_config of ANDgate5 is
   for untitled
   end for;
end ANDgate5_config;