configuration ANDgate_config of ANDgate is
   for untitled
   end for;
end ANDgate_config;