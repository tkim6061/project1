configuration ORgate3_config of ORgate3 is
   for untitled
   end for;
end ORgate3_config;