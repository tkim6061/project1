configuration ORgate4_config of ORgate4 is
   for untitled
   end for;
end ORgate4_config;