-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
configuration scrambler_config of scrambler is
   for struct
   end for;
end scrambler_config;
