-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
configuration Corrector_config of Corrector is
   for struct
   end for;
end Corrector_config;
