configuration ANDgate3_config of ANDgate3 is
   for untitled
   end for;
end ANDgate3_config;