configuration ORgate5_config of ORgate5 is
   for untitled
   end for;
end ORgate5_config;