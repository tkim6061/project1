configuration XORgate_config of XORgate is
   for untitled
   end for;
end XORgate_config;